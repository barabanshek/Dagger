// Author: Cornell University
//
// Module Name :    nic_defs
// Project :        F-NIC
// Description :    Definitions for the NIC module
//

`ifndef NIC_DEFS_VH_
`define NIC_DEFS_VH_

`include "cpu_if_defs.vh"

parameter LMAX_CCIP_BATCH = 2;
parameter LMAX_CCIP_DMA_BATCH = 6;

// RPC interfaces
typedef struct packed {
    logic [7:0] flow_id;    //TODO: it's a temporary solution, will have an RPC descriptor table later
    RpcPckt     rpc_data;
} RpcIf;

// Network interfaces
localparam TRANSPORT_DATA_WIDTH = 512;

typedef struct packed {
    logic[31:0]             payload_size;
    logic[31:0]             conn_id;
} NetworkPacketHdr;

typedef struct packed {
    NetworkPacketHdr hdr;
    logic[TRANSPORT_DATA_WIDTH-1:0] payload;
} NetworkPacketInternal;


`endif //  NIC_DEFS_VH_
